module Counter_divider(
	//entrada de dados
	clk,
	
	//saída de dados
	clk1,
	clk2,
	clk3,
	clk4
);

	// Input Port(s)
	input wire clk;
	
	// Output Port(s)
	output wire clk1;  //wire ou reg?
	output wire clk2;  //wire ou reg?
	output wire clk3;  //wire ou reg?
	output wire clk4;  //wire ou reg?
endmodule