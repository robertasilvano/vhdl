module Counter_divider(
clk,
clk1,
clk2,
clk3,
clk4
);

	input wire clk;
	input wire clk1;
	input wire clk2;
	input wire clk3;
	input wire clk4;
endmodule