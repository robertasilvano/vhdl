library verilog;
use verilog.vl_types.all;
entity Topo_tb is
end Topo_tb;
