module Dec7seg(
G,
O
);

	localparam p_G = 4;
	localparam p_O = 7;

	input wire [p_G - 1:0] G;
	input wire [p_O - 1:0] O;
endmodule
